--  Copyright 2020 Equinor ASA
--
--  This file is part of the Open Porous Media project (OPM).
--
--  OPM is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  OPM is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with OPM.  If not, see <http://www.gnu.org/licenses/>.

-- ******************************
-- top for AXI memory read module
-- ******************************
-- WARNING: this design is meant for a read port connected to DDR memory.
-- This design integrates:
-- * the read_input core generated by HLS
-- * the AXI master core generated by HLS
-- * a FIFO that includes the almost_empty signal, with separate clock domains
-- * registers for address, data_len, offset when ap_start is set (HLS
--   module does not properly register them!)

-- FIXME: these signals can be considered as static when they cross clock domains,
-- but a timing exception must be applied to them:
--   address_r, data_len_r, mem_offset_r

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
library xpm;
  use xpm.vcomponents.all;
library work;
  use work.axi_io_common.all;
  use work.constants.all;

entity mem_read_top_async_ddr is
port (
  -- HLS/parameters interface
  clk_rd : in std_logic;
  rst_rd : in std_logic;
  ap_start : in std_logic;
  ap_done : out std_logic;
  ap_idle : out std_logic;
  ap_ready : out std_logic;
  fifo_busy : out std_logic;
  address : in std_logic_vector (63 downto 0);
  data_len : in std_logic_vector (31 downto 0);
  mem_offset : in std_logic_vector (63 downto 0);
  -- FIFO (stream) interface - uses clk_rd
  in_fifo_data : out std_logic_vector(C_FIFOREAD_DATAOUT_WIDTH-1 downto 0);
  in_fifo_empty : out std_logic;
  in_fifo_almost_empty : out std_logic;
  in_fifo_rd : in std_logic;
  -- AXI interface
  clk_axi : in std_logic;
  rst_axi : in std_logic;
  m_axi_gmem_AWVALID : out std_logic;
  m_axi_gmem_AWREADY : in std_logic;
  m_axi_gmem_AWADDR : out std_logic_vector (C_M_AXI_GMEMREAD_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_AWID : out std_logic_vector (C_M_AXI_GMEMREAD_ID_WIDTH-1 downto 0);
  m_axi_gmem_AWLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_AWSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWUSER : out std_logic_vector (C_M_AXI_GMEMREAD_AWUSER_WIDTH-1 downto 0);
  m_axi_gmem_WVALID : out std_logic;
  m_axi_gmem_WREADY : in std_logic;
  m_axi_gmem_WDATA : out std_logic_vector (C_M_AXI_GMEMREAD_DATA_WIDTH-1 downto 0);
  m_axi_gmem_WSTRB : out std_logic_vector (C_M_AXI_GMEMREAD_DATA_WIDTH/8-1 downto 0);
  m_axi_gmem_WLAST : out std_logic;
  m_axi_gmem_WID : out std_logic_vector (C_M_AXI_GMEMREAD_ID_WIDTH-1 downto 0);
  m_axi_gmem_WUSER : out std_logic_vector (C_M_AXI_GMEMREAD_WUSER_WIDTH-1 downto 0);
  m_axi_gmem_ARVALID : out std_logic;
  m_axi_gmem_ARREADY : in std_logic;
  m_axi_gmem_ARADDR : out std_logic_vector (C_M_AXI_GMEMREAD_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_ARID : out std_logic_vector (C_M_AXI_GMEMREAD_ID_WIDTH-1 downto 0);
  m_axi_gmem_ARLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_ARSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARUSER : out std_logic_vector (C_M_AXI_GMEMREAD_ARUSER_WIDTH-1 downto 0);
  m_axi_gmem_RVALID : in std_logic;
  m_axi_gmem_RREADY : out std_logic;
  m_axi_gmem_RDATA : in std_logic_vector (C_M_AXI_GMEMREAD_DATA_WIDTH-1 downto 0);
  m_axi_gmem_RLAST : in std_logic;
  m_axi_gmem_RID : in std_logic_vector (C_M_AXI_GMEMREAD_ID_WIDTH-1 downto 0);
  m_axi_gmem_RUSER : in std_logic_vector (C_M_AXI_GMEMREAD_RUSER_WIDTH-1 downto 0);
  m_axi_gmem_RRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BVALID : in std_logic;
  m_axi_gmem_BREADY : out std_logic;
  m_axi_gmem_BRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BID : in std_logic_vector (C_M_AXI_GMEMREAD_ID_WIDTH-1 downto 0);
  m_axi_gmem_BUSER : in std_logic_vector (C_M_AXI_GMEMREAD_BUSER_WIDTH-1 downto 0)
);
end;

architecture behavioral of mem_read_top_async_ddr is
signal axi_ap_start, axi_ap_done, axi_ap_idle, axi_ap_ready: std_logic;
signal reg_ap_start, reg_ap_done, reg_ap_idle, reg_ap_ready: std_logic;
signal fifo_wr_busy, fifo_wr_busy_clkrd, fifo_rd_busy: std_logic;
signal address_r,reg_address: std_logic_vector (63 downto 0);
signal data_len_r,reg_data_len: std_logic_vector (31 downto 0);
signal mem_offset_r: std_logic_vector(63 downto 0);
signal reg_mem_offset_shifted: std_logic_vector(57 downto 0);
signal read_input_fifo_data: std_logic_vector(C_FIFOREAD_DATAIN_WIDTH-1 downto 0);
signal read_input_fifo_full_n, read_input_fifo_wr: std_logic;
signal read_input_m_axi_in_V_ARVALID: std_logic;
signal read_input_m_axi_in_V_ARREADY: std_logic;
signal read_input_m_axi_in_V_ARADDR: std_logic_vector (63 downto 0);
signal read_input_m_axi_in_V_ARID: std_logic_vector (0 downto 0);
signal read_input_m_axi_in_V_ARLEN: std_logic_vector (31 downto 0);
signal read_input_m_axi_in_V_ARSIZE: std_logic_vector (2 downto 0);
signal read_input_m_axi_in_V_ARLOCK: std_logic_vector (1 downto 0);
signal read_input_m_axi_in_V_ARCACHE: std_logic_vector (3 downto 0);
signal read_input_m_axi_in_V_ARQOS: std_logic_vector (3 downto 0);
signal read_input_m_axi_in_V_ARPROT: std_logic_vector (2 downto 0);
signal read_input_m_axi_in_V_ARUSER: std_logic_vector (0 downto 0);
signal read_input_m_axi_in_V_ARBURST: std_logic_vector (1 downto 0);
signal read_input_m_axi_in_V_ARREGION: std_logic_vector (3 downto 0);
signal read_input_m_axi_in_V_RVALID: std_logic;
signal read_input_m_axi_in_V_RREADY: std_logic;
signal read_input_m_axi_in_V_RDATA: std_logic_vector (511 downto 0);
signal read_input_m_axi_in_V_RID: std_logic_vector (0 downto 0);
signal read_input_m_axi_in_V_RUSER: std_logic_vector (0 downto 0);
signal read_input_m_axi_in_V_RRESP: std_logic_vector (1 downto 0);
signal read_input_m_axi_in_V_RLAST: std_logic;
type control_t is (idle,running);
-- number of words contained by the FIFO
constant FIFO_WORDS: integer := 512;

begin

--******************************************************************************
-- clock domain: clk_rd
--******************************************************************************

  -- register address, data_len, mem_offset in clk_rd domain when ap_start is
  -- set (there is no guarantee they'll be valid afterwards)
  control_start_p: process(clk_rd)
  begin
    if rising_edge(clk_rd) then
      if rst_rd = '1' then
        address_r <= (others => '0');
        data_len_r <= (others => '0');
        mem_offset_r <= (others => '0');
      elsif (ap_start = '1') then
        address_r <= address;
        data_len_r <= data_len;
        mem_offset_r <= mem_offset;
      end if;
    end if;
  end process;

  -- fifo_busy signal is a summary of if_wr_busy and if_rd_busy, syncronized to clk_rd
  fifo_busy <= fifo_wr_busy_clkrd or fifo_rd_busy;

--******************************************************************************
-- clock domain: BOTH
--******************************************************************************

  -- read data FIFO
  indata_fifo_i: entity work.fifo_in_async_w512
  generic map (
    MEM_STYLE  => "block",
    DATA_WIDTH => 512,
    DEPTH      => FIFO_WORDS)
  port map (
    reset => rst_axi,
    clk_wr => clk_axi,
    if_wr_busy => fifo_wr_busy,
    if_write => read_input_fifo_wr,
    if_din => read_input_fifo_data,
    if_almost_full => open,
    if_full_n => read_input_fifo_full_n,
    clk_rd => clk_rd,
    if_rd_busy => fifo_rd_busy,
    if_read => in_fifo_rd,
    if_dout => in_fifo_data,
    if_almost_empty => in_fifo_almost_empty,
    if_empty => in_fifo_empty
  );

--******************************************************************************
-- CDC logic
--******************************************************************************

  -- CDC for HLS interface - pulse signal ap_start
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_start_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => 4,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_rd,
    src_rst => '0', --rst_rd,
    src_pulse => ap_start, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_axi,
    dest_rst => '0', --rst_axi,
    dest_pulse =>  axi_ap_start -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - pulse signal ap_done
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_done_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => 4,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_axi,
    src_rst => '0', --rst_axi,
    src_pulse => axi_ap_done, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_rd,
    dest_rst => '0', --rst_rd,
    dest_pulse =>  ap_done -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - pulse signal ap_ready
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_ready_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => 4,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_axi,
    src_rst => '0', --rst_axi,
    src_pulse => axi_ap_ready, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_rd,
    dest_rst => '0', --rst_rd,
    dest_pulse =>  ap_ready -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - non-pulse signal ap_idle
  -- xpm_cdc_single: Single-bit Synchronizer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_idle_cdc_i: xpm_cdc_single
  generic map (
    DEST_SYNC_FF => 4,   -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 0,   -- 0=disable simulation init values, 1=enable simulation init values
    SIM_ASSERT_CHK => 1, -- 0=disable simulation messages, 1=enable simulation messages
    SRC_INPUT_REG => 1   -- 0=do not register input, 1=register input
  )
  port map (
    src_clk => clk_axi,  -- optional; required when SRC_INPUT_REG = 1
    src_in => axi_ap_idle,
    dest_clk => clk_rd,
    dest_out => ap_idle
  );

  -- CDC for non-pulse signal if_wr_busy
  -- xpm_cdc_single: Single-bit Synchronizer
  -- Xilinx Parameterized Macro, version 2019.2
  if_wr_busy_cdc_i: xpm_cdc_single
  generic map (
    DEST_SYNC_FF => 4,   -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 0,   -- 0=disable simulation init values, 1=enable simulation init values
    SIM_ASSERT_CHK => 1, -- 0=disable simulation messages, 1=enable simulation messages
    SRC_INPUT_REG => 1   -- 0=do not register input, 1=register input
  )
  port map (
    src_clk => clk_axi,  -- optional; required when SRC_INPUT_REG = 1
    src_in => fifo_wr_busy,
    dest_clk => clk_rd,
    dest_out => fifo_wr_busy_clkrd
  );

--******************************************************************************
-- clock domain: clk_axi
--******************************************************************************

  -- process to resync the signals that must be registered to fix the wrong
  -- bevahior of read_input unit
  -- uses single-shot style for axi_ap_done
  control_os_p: process(clk_axi, axi_ap_start)
  variable state: control_t;
  variable vready: std_logic;
  begin
    if rising_edge(clk_axi) then
      if rst_axi = '1' then
        axi_ap_done <= '0';
        axi_ap_ready <= '0';
        vready := '0';
        reg_ap_start <= '0';
        state := idle;
      else
        case state is
          when idle =>
            -- wait until axi_ap_start is set
            axi_ap_done <= '0';
            axi_ap_ready <= '0';
            vready := '0';
            reg_ap_start <= '0';
            if (axi_ap_start = '1') then
              reg_ap_start <= '1';
              reg_address <= address_r;
              reg_data_len <= data_len_r;
              reg_mem_offset_shifted <= mem_offset_r(63 downto 6);
              state := running;
            end if;
          when running =>
            -- run the unit
            reg_ap_start <= '0';
            if (reg_ap_done = '1') then
              axi_ap_done <= '1';
              axi_ap_ready <= '1';
              vready := '1';
              state := idle;
            end if;
          when others =>
            state := idle;
        end case;
      end if;
    end if;
    if (axi_ap_start = '1') or (vready = '1') or (state = running) then
      axi_ap_idle <= '0';
    else
      axi_ap_idle <= '1';
    end if;
  end process;

  -- memory read module
  read_input_i: entity work.read_input
  port map (
    ap_clk => clk_axi,
    ap_rst => rst_axi,
    ap_start => reg_ap_start,
    ap_done => reg_ap_done,
    ap_idle => reg_ap_idle,
    ap_ready => reg_ap_ready,
    m_axi_in_V_AWVALID => open,
    m_axi_in_V_AWREADY => '0',
    m_axi_in_V_AWADDR => open,
    m_axi_in_V_AWID => open,
    m_axi_in_V_AWLEN => open,
    m_axi_in_V_AWSIZE => open,
    m_axi_in_V_AWBURST => open,
    m_axi_in_V_AWLOCK => open,
    m_axi_in_V_AWCACHE => open,
    m_axi_in_V_AWPROT => open,
    m_axi_in_V_AWQOS => open,
    m_axi_in_V_AWREGION => open,
    m_axi_in_V_AWUSER => open,
    m_axi_in_V_WVALID => open,
    m_axi_in_V_WREADY => '0',
    m_axi_in_V_WDATA => open,
    m_axi_in_V_WSTRB => open,
    m_axi_in_V_WLAST => open,
    m_axi_in_V_WID => open,
    m_axi_in_V_WUSER => open,
    m_axi_in_V_ARVALID => read_input_m_axi_in_V_ARVALID,
    m_axi_in_V_ARREADY => read_input_m_axi_in_V_ARREADY,
    m_axi_in_V_ARADDR => read_input_m_axi_in_V_ARADDR,
    m_axi_in_V_ARID => read_input_m_axi_in_V_ARID,
    m_axi_in_V_ARLEN => read_input_m_axi_in_V_ARLEN,
    m_axi_in_V_ARSIZE => read_input_m_axi_in_V_ARSIZE,
    m_axi_in_V_ARBURST => read_input_m_axi_in_V_ARBURST,
    m_axi_in_V_ARLOCK => read_input_m_axi_in_V_ARLOCK,
    m_axi_in_V_ARCACHE => read_input_m_axi_in_V_ARCACHE,
    m_axi_in_V_ARPROT => read_input_m_axi_in_V_ARPROT,
    m_axi_in_V_ARQOS => read_input_m_axi_in_V_ARQOS,
    m_axi_in_V_ARREGION => read_input_m_axi_in_V_ARREGION,
    m_axi_in_V_ARUSER => read_input_m_axi_in_V_ARUSER,
    m_axi_in_V_RVALID => read_input_m_axi_in_V_RVALID,
    m_axi_in_V_RREADY => read_input_m_axi_in_V_RREADY,
    m_axi_in_V_RDATA => read_input_m_axi_in_V_RDATA,
    m_axi_in_V_RLAST => read_input_m_axi_in_V_RLAST,
    m_axi_in_V_RID => read_input_m_axi_in_V_RID,
    m_axi_in_V_RUSER => read_input_m_axi_in_V_RUSER,
    m_axi_in_V_RRESP => read_input_m_axi_in_V_RRESP,
    m_axi_in_V_BVALID => '0',
    m_axi_in_V_BREADY => open,
    m_axi_in_V_BRESP => "00",
    m_axi_in_V_BID => "0",
    m_axi_in_V_BUSER => "0",
    in_V_offset => reg_mem_offset_shifted,
    address => reg_address,
    data_len => reg_data_len,
    elemStream_V_V_din => read_input_fifo_data,
    elemStream_V_V_full_n => read_input_fifo_full_n,
    elemStream_V_V_write => read_input_fifo_wr
  );

  -- AXI interface
  hls_m_axi_i: entity work.hls_sdaccel_kernel_iostreams_hls_gmem0_m_axi
  generic map (
    CONSERVATIVE => 0,
    USER_DW => 512,
    USER_AW => 64,
    USER_MAXREQS => 8,           -- do not set below 2
    NUM_READ_OUTSTANDING => 8,   -- do not set below 2
    NUM_WRITE_OUTSTANDING => 2,  -- do not set below 2 - no writes in this module
    MAX_READ_BURST_LENGTH => 256,
    MAX_WRITE_BURST_LENGTH => 2, -- no writes in this module
    C_M_AXI_ID_WIDTH => C_M_AXI_GMEMREAD_ID_WIDTH,
    C_M_AXI_ADDR_WIDTH => C_M_AXI_GMEMREAD_ADDR_WIDTH,
    C_TARGET_ADDR => 16#00000000#,
    C_M_AXI_DATA_WIDTH => C_M_AXI_GMEMREAD_DATA_WIDTH,
    C_M_AXI_AWUSER_WIDTH => C_M_AXI_GMEMREAD_AWUSER_WIDTH,
    C_M_AXI_ARUSER_WIDTH => C_M_AXI_GMEMREAD_ARUSER_WIDTH,
    C_M_AXI_WUSER_WIDTH => C_M_AXI_GMEMREAD_WUSER_WIDTH,
    C_M_AXI_RUSER_WIDTH => C_M_AXI_GMEMREAD_RUSER_WIDTH,
    C_M_AXI_BUSER_WIDTH => C_M_AXI_GMEMREAD_BUSER_WIDTH,
    C_USER_VALUE => C_M_AXI_GMEMREAD_USER_VALUE,
    C_PROT_VALUE => C_M_AXI_GMEMREAD_PROT_VALUE,
    C_CACHE_VALUE => C_M_AXI_GMEMREAD_CACHE_VALUE)
  port map (
    ACLK => clk_axi,
    ARESET => rst_axi,
    ACLK_EN => '1',
    AWVALID => m_axi_gmem_AWVALID,
    AWREADY => m_axi_gmem_AWREADY,
    AWADDR => m_axi_gmem_AWADDR,
    AWID => m_axi_gmem_AWID,
    AWLEN => m_axi_gmem_AWLEN,
    AWSIZE => m_axi_gmem_AWSIZE,
    AWBURST => m_axi_gmem_AWBURST,
    AWLOCK => m_axi_gmem_AWLOCK,
    AWCACHE => m_axi_gmem_AWCACHE,
    AWPROT => m_axi_gmem_AWPROT,
    AWQOS => m_axi_gmem_AWQOS,
    AWREGION => m_axi_gmem_AWREGION,
    AWUSER => m_axi_gmem_AWUSER,
    WVALID => m_axi_gmem_WVALID,
    WREADY => m_axi_gmem_WREADY,
    WDATA => m_axi_gmem_WDATA,
    WSTRB => m_axi_gmem_WSTRB,
    WLAST => m_axi_gmem_WLAST,
    WID => m_axi_gmem_WID,
    WUSER => m_axi_gmem_WUSER,
    ARVALID => m_axi_gmem_ARVALID,
    ARREADY => m_axi_gmem_ARREADY,
    ARADDR => m_axi_gmem_ARADDR,
    ARID => m_axi_gmem_ARID,
    ARLEN => m_axi_gmem_ARLEN,
    ARSIZE => m_axi_gmem_ARSIZE,
    ARBURST => m_axi_gmem_ARBURST,
    ARLOCK => m_axi_gmem_ARLOCK,
    ARCACHE => m_axi_gmem_ARCACHE,
    ARPROT => m_axi_gmem_ARPROT,
    ARQOS => m_axi_gmem_ARQOS,
    ARREGION => m_axi_gmem_ARREGION,
    ARUSER => m_axi_gmem_ARUSER,
    RVALID => m_axi_gmem_RVALID,
    RREADY => m_axi_gmem_RREADY,
    RDATA => m_axi_gmem_RDATA,
    RLAST => m_axi_gmem_RLAST,
    RID => m_axi_gmem_RID,
    RUSER => m_axi_gmem_RUSER,
    RRESP => m_axi_gmem_RRESP,
    BVALID => m_axi_gmem_BVALID,
    BREADY => m_axi_gmem_BREADY,
    BRESP => m_axi_gmem_BRESP,
    BID => m_axi_gmem_BID,
    BUSER => m_axi_gmem_BUSER,
    -- internal bus ports
    -- write channel is disabled for this module
    I_AWVALID => '0',
    I_AWREADY => open,
    I_AWADDR => x"0000000000000000",
    I_AWID => "0",
    I_AWLEN => x"00000000",
    I_AWSIZE => "000",
    I_AWLOCK => "00",
    I_AWCACHE => "0000",
    I_AWQOS => "0000",
    I_AWPROT => "000",
    I_AWUSER => "0",
    I_AWBURST => "00",
    I_AWREGION => "0000",
    I_WVALID => '0',
    I_WREADY => open,
    I_WDATA => ap_const_lv512_lc_1,
    I_WID => "0",
    I_WUSER => "0",
    I_WLAST => '0',
    I_WSTRB => x"0000000000000000",
    I_ARVALID => read_input_m_axi_in_V_ARVALID,
    I_ARREADY => read_input_m_axi_in_V_ARREADY,
    I_ARADDR => read_input_m_axi_in_V_ARADDR,
    I_ARID => read_input_m_axi_in_V_ARID,
    I_ARLEN => read_input_m_axi_in_V_ARLEN,
    I_ARSIZE => read_input_m_axi_in_V_ARSIZE,
    I_ARLOCK => read_input_m_axi_in_V_ARLOCK,
    I_ARCACHE => read_input_m_axi_in_V_ARCACHE,
    I_ARQOS => read_input_m_axi_in_V_ARQOS,
    I_ARPROT => read_input_m_axi_in_V_ARPROT,
    I_ARUSER => read_input_m_axi_in_V_ARUSER,
    I_ARBURST => read_input_m_axi_in_V_ARBURST,
    I_ARREGION => read_input_m_axi_in_V_ARREGION,
    I_RVALID => read_input_m_axi_in_V_RVALID,
    I_RREADY => read_input_m_axi_in_V_RREADY,
    I_RDATA => read_input_m_axi_in_V_RDATA,
    I_RID => read_input_m_axi_in_V_RID,
    I_RUSER => read_input_m_axi_in_V_RUSER,
    I_RRESP => read_input_m_axi_in_V_RRESP,
    I_RLAST => read_input_m_axi_in_V_RLAST,
    I_BVALID => open,
    I_BREADY => '0',
    I_BRESP => open,
    I_BID => open,
    I_BUSER => open
  );

end architecture;

