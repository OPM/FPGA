../output-impl-vhdl/write_output_buffer_V.vhd