../output-impl-vhdl/read_memory_proc.vhd