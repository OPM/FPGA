--  Copyright 2020 Equinor ASA
--
--  This file is part of the Open Porous Media project (OPM).
--
--  OPM is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  OPM is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with OPM.  If not, see <http://www.gnu.org/licenses/>.

-- *******************************
-- top for AXI memory write module
-- *******************************
-- WARNING: this design is meant for a write port connected to HBM memory.
-- This design integrates:
-- * the write_output core generated by HLS
-- * the AXI master core generated by HLS
-- * a FIFO that includes the almost_full signal (generated by HLS and modified)
-- * registers for address, data_len, offset when ap_start is set (HLS
--   module does not properly register them!)

-- FIXME: these signals can be considered as static when they cross clock domains,
-- but a timing exception must be applied to them:
--   address_r, data_len_r, mem_offset_r

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
library xpm;
  use xpm.vcomponents.all;
library work;
  use work.axi_io_common.all;
  use work.constants.all;

entity mem_write_top_async_hbm is
port (
  -- HLS/parameters interface
  clk_wr : in std_logic;
  rst_wr : in std_logic;
  ap_start : in std_logic;
  ap_done : out std_logic;
  ap_idle : out std_logic;
  ap_ready : out std_logic;
  fifo_busy : out std_logic;
  address : in std_logic_vector (63 downto 0);
  data_len : in std_logic_vector (31 downto 0);
  mem_offset : in std_logic_vector (63 downto 0);
  -- FIFO (stream) interface - uses clk_wr
  out_fifo_data : in std_logic_vector(C_FIFOWRITE_DATAIN_WIDTH-1 downto 0);
  out_fifo_full : out std_logic;
  out_fifo_almost_full : out std_logic;
  out_fifo_wr : in std_logic;
  -- AXI interface
  clk_axi : in std_logic;
  rst_axi : in std_logic;
  m_axi_gmem_AWVALID : out std_logic;
  m_axi_gmem_AWREADY : in std_logic;
  m_axi_gmem_AWADDR : out std_logic_vector (C_M_AXI_GMEMWRITE_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_AWID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_AWLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_AWSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_AWUSER_WIDTH-1 downto 0);
  m_axi_gmem_WVALID : out std_logic;
  m_axi_gmem_WREADY : in std_logic;
  m_axi_gmem_WDATA : out std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH-1 downto 0);
  m_axi_gmem_WSTRB : out std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH/8-1 downto 0);
  m_axi_gmem_WLAST : out std_logic;
  m_axi_gmem_WID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_WUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_WUSER_WIDTH-1 downto 0);
  m_axi_gmem_ARVALID : out std_logic;
  m_axi_gmem_ARREADY : in std_logic;
  m_axi_gmem_ARADDR : out std_logic_vector (C_M_AXI_GMEMWRITE_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_ARID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_ARLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_ARSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_ARUSER_WIDTH-1 downto 0);
  m_axi_gmem_RVALID : in std_logic;
  m_axi_gmem_RREADY : out std_logic;
  m_axi_gmem_RDATA : in std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH-1 downto 0);
  m_axi_gmem_RLAST : in std_logic;
  m_axi_gmem_RID : in std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_RUSER : in std_logic_vector (C_M_AXI_GMEMWRITE_RUSER_WIDTH-1 downto 0);
  m_axi_gmem_RRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BVALID : in std_logic;
  m_axi_gmem_BREADY : out std_logic;
  m_axi_gmem_BRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BID : in std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_BUSER : in std_logic_vector (C_M_AXI_GMEMWRITE_BUSER_WIDTH-1 downto 0)
);
end;

architecture behavioral of mem_write_top_async_hbm is
signal axi_ap_start, axi_ap_done, axi_ap_idle, axi_ap_ready: std_logic;
signal reg_ap_start, reg_ap_done, reg_ap_idle, reg_ap_ready: std_logic;
signal fifo_wr_busy, fifo_rd_busy, fifo_rd_busy_clkwr: std_logic;
signal address_r,reg_address: std_logic_vector (63 downto 0);
signal data_len_r,reg_data_len: std_logic_vector (31 downto 0);
signal mem_offset_r: std_logic_vector(63 downto 0);
-- keep the registered parameter signals as they will be used to specify a timing exception
attribute dont_touch: string;
attribute dont_touch of address_r: signal is "true";
attribute dont_touch of data_len_r: signal is "true";
attribute dont_touch of mem_offset_r: signal is "true";
signal reg_mem_offset_shifted: std_logic_vector(57 downto 0);
signal write_output_fifo_data: std_logic_vector(C_FIFOWRITE_DATAOUT_WIDTH-1 downto 0);
signal write_output_fifo_empty_n, write_output_fifo_rd: std_logic;
signal write_output_m_axi_out_V_AWVALID: std_logic;
signal write_output_m_axi_out_V_AWREADY: std_logic;
signal write_output_m_axi_out_V_AWADDR: std_logic_vector (63 downto 0);
signal write_output_m_axi_out_V_AWID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_AWLEN: std_logic_vector (31 downto 0);
signal write_output_m_axi_out_V_AWSIZE: std_logic_vector (2 downto 0);
signal write_output_m_axi_out_V_AWLOCK: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_AWCACHE: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_AWQOS: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_AWPROT: std_logic_vector (2 downto 0);
signal write_output_m_axi_out_V_AWUSER: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_AWBURST: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_AWREGION: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_WVALID: std_logic;
signal write_output_m_axi_out_V_WREADY: std_logic;
signal write_output_m_axi_out_V_WDATA: std_logic_vector (511 downto 0);
signal write_output_m_axi_out_V_WID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_WUSER: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_WLAST: std_logic;
signal write_output_m_axi_out_V_WSTRB: std_logic_vector (63 downto 0);
signal write_output_m_axi_out_V_BVALID: std_logic;
signal write_output_m_axi_out_V_BREADY: std_logic;
signal write_output_m_axi_out_V_BRESP: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_BID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_BUSER: std_logic_vector (0 downto 0);
type control_t is (idle,running);
-- number of words contained by the FIFO
constant FIFO_WORDS: integer := 256;

begin

--******************************************************************************
-- clock domain: clk_wr
--******************************************************************************

  -- register address, data_len, mem_offset in clk_wr domain when ap_start is
  -- set (there is no guarantee they'll be valid afterwards)
  control_start_p: process(clk_wr)
  begin
    if rising_edge(clk_wr) then
      if rst_wr = '1' then
        address_r <= (others => '0');
        data_len_r <= (others => '0');
        mem_offset_r <= (others => '0');
      elsif (ap_start = '1') then
        address_r <= address;
        data_len_r <= data_len;
        mem_offset_r <= mem_offset;
      end if;
    end if;
  end process;

  -- fifo_busy signal is a summary of if_wr_busy and if_rd_busy, syncronized to clk_wr
  fifo_busy <= fifo_wr_busy or fifo_rd_busy_clkwr;

--******************************************************************************
-- clock domain: BOTH
--******************************************************************************

  -- write data FIFO
  outdata_fifo_i: entity work.fifo_out_async_w512
  generic map (
    MEM_STYLE  => "block",
    DATA_WIDTH => 512,
    DEPTH      => FIFO_WORDS)
  port map (
    reset => rst_wr,
    clk_wr => clk_wr,
    if_wr_busy => fifo_wr_busy,
    if_write => out_fifo_wr,
    if_din => out_fifo_data,
    if_almost_full => out_fifo_almost_full,
    if_full => out_fifo_full,
    clk_rd => clk_axi,
    if_rd_busy => fifo_rd_busy,
    if_read => write_output_fifo_rd,
    if_dout => write_output_fifo_data,
    if_almost_empty => open,
    if_empty_n => write_output_fifo_empty_n
  );

--******************************************************************************
-- CDC logic
--******************************************************************************

  -- CDC for HLS interface - pulse signal ap_start
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_start_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => CDC_STAGES_PULSE,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_wr,
    src_rst => '0', --rst_wr,
    src_pulse => ap_start, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_axi,
    dest_rst => '0', --rst_axi,
    dest_pulse =>  axi_ap_start -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - pulse signal ap_done
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_done_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => CDC_STAGES_PULSE,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_axi,
    src_rst => '0', --rst_axi,
    src_pulse => axi_ap_done, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_wr,
    dest_rst => '0', --rst_wr,
    dest_pulse =>  ap_done -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - pulse signal ap_ready
  -- xpm_cdc_pulse: Pulse Transfer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_ready_cdc_i: xpm_cdc_pulse
  generic map (
    DEST_SYNC_FF => CDC_STAGES_PULSE,  -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 1,  -- 0=disable simulation init values, 1=enable simulation init values
    REG_OUTPUT => 1,    -- 0=disable registered output, 1=enable registered output
    RST_USED => 0,      -- 0=no reset, 1=implement reset
    SIM_ASSERT_CHK => 1 -- 0=disable simulation messages, 1=enable simulation messages
  )
  port map (
    src_clk => clk_axi,
    src_rst => '0', --rst_axi,
    src_pulse => axi_ap_ready, -- Min gap between pulses must be 2*(larger(src_clk period, dest_clk period))
    dest_clk => clk_wr,
    dest_rst => '0', --rst_wr,
    dest_pulse =>  ap_ready -- This output is combinatorial unless REG_OUTPUT is set to 1.
  );

  -- CDC for HLS interface - non-pulse signal ap_idle
  -- xpm_cdc_single: Single-bit Synchronizer
  -- Xilinx Parameterized Macro, version 2019.2
  ap_idle_cdc_i: xpm_cdc_single
  generic map (
    DEST_SYNC_FF => CDC_STAGES_SINGLE,   -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 0,   -- 0=disable simulation init values, 1=enable simulation init values
    SIM_ASSERT_CHK => 1, -- 0=disable simulation messages, 1=enable simulation messages
    SRC_INPUT_REG => 1   -- 0=do not register input, 1=register input
  )
  port map (
    src_clk => clk_axi,  -- optional; required when SRC_INPUT_REG = 1
    src_in => axi_ap_idle,
    dest_clk => clk_wr,
    dest_out => ap_idle
  );

  -- CDC for non-pulse signal if_rd_busy
  -- xpm_cdc_single: Single-bit Synchronizer
  -- Xilinx Parameterized Macro, version 2019.2
  if_rd_busy_cdc_i: xpm_cdc_single
  generic map (
    DEST_SYNC_FF => CDC_STAGES_SINGLE,   -- Number of register stages; range: 2-10
    INIT_SYNC_FF => 0,   -- 0=disable simulation init values, 1=enable simulation init values
    SIM_ASSERT_CHK => 1, -- 0=disable simulation messages, 1=enable simulation messages
    SRC_INPUT_REG => 1   -- 0=do not register input, 1=register input
  )
  port map (
    src_clk => clk_axi,  -- optional; required when SRC_INPUT_REG = 1
    src_in => fifo_rd_busy,
    dest_clk => clk_wr,
    dest_out => fifo_rd_busy_clkwr
  );

--******************************************************************************
-- clock domain: clk_axi
--******************************************************************************

  -- process to resync the signals that must be registered to fix the wrong
  -- bevahior of write_output unit
  -- uses single-shot style for axi_ap_done
  control_os_p: process(clk_axi, axi_ap_start)
  variable state: control_t;
  variable vready: std_logic;
  begin
    if rising_edge(clk_axi) then
      if rst_axi = '1' then
        axi_ap_done <= '0';
        axi_ap_ready <= '0';
        vready := '0';
        reg_ap_start <= '0';
        state := idle;
      else
        case state is
          when idle =>
            -- wait until ap_start is set
            axi_ap_done <= '0';
            axi_ap_ready <= '0';
            vready := '0';
            reg_ap_start <= '0';
            if (axi_ap_start = '1') then
              reg_ap_start <= '1';
              reg_address <= address_r;
              reg_data_len <= data_len_r;
              reg_mem_offset_shifted <= mem_offset_r(63 downto 6);
              state := running;
            end if;
          when running =>
            -- run the unit
            reg_ap_start <= '0';
            if (reg_ap_done = '1') then
              axi_ap_done <= '1';
              axi_ap_ready <= '1';
              vready := '1';
              state := idle;
            end if;
          when others =>
            state := idle;
        end case;
      end if;
    end if;
    if (axi_ap_start = '1') or (vready = '1') or (state = running) then
      axi_ap_idle <= '0';
    else
      axi_ap_idle <= '1';
    end if;
  end process;

  -- memory write module
  write_output_i: entity work.write_output
  port map (
    ap_clk => clk_axi,
    ap_rst => rst_axi,
    ap_start => reg_ap_start,
    ap_done => reg_ap_done,
    ap_idle => reg_ap_idle,
    ap_ready => reg_ap_ready,
    resultStream_V_V_dout => write_output_fifo_data,
    resultStream_V_V_empty_n => write_output_fifo_empty_n,
    resultStream_V_V_read => write_output_fifo_rd,
    m_axi_out_V_AWVALID => write_output_m_axi_out_V_AWVALID,
    m_axi_out_V_AWREADY => write_output_m_axi_out_V_AWREADY,
    m_axi_out_V_AWADDR => write_output_m_axi_out_V_AWADDR,
    m_axi_out_V_AWID => write_output_m_axi_out_V_AWID,
    m_axi_out_V_AWLEN => write_output_m_axi_out_V_AWLEN,
    m_axi_out_V_AWSIZE => write_output_m_axi_out_V_AWSIZE,
    m_axi_out_V_AWBURST => write_output_m_axi_out_V_AWBURST,
    m_axi_out_V_AWLOCK => write_output_m_axi_out_V_AWLOCK,
    m_axi_out_V_AWCACHE => write_output_m_axi_out_V_AWCACHE,
    m_axi_out_V_AWPROT => write_output_m_axi_out_V_AWPROT,
    m_axi_out_V_AWQOS => write_output_m_axi_out_V_AWQOS,
    m_axi_out_V_AWREGION => write_output_m_axi_out_V_AWREGION,
    m_axi_out_V_AWUSER => write_output_m_axi_out_V_AWUSER,
    m_axi_out_V_WVALID => write_output_m_axi_out_V_WVALID,
    m_axi_out_V_WREADY => write_output_m_axi_out_V_WREADY,
    m_axi_out_V_WDATA => write_output_m_axi_out_V_WDATA,
    m_axi_out_V_WSTRB => write_output_m_axi_out_V_WSTRB,
    m_axi_out_V_WLAST => write_output_m_axi_out_V_WLAST,
    m_axi_out_V_WID => write_output_m_axi_out_V_WID,
    m_axi_out_V_WUSER => write_output_m_axi_out_V_WUSER,
    m_axi_out_V_ARVALID => open,
    m_axi_out_V_ARREADY => '0',
    m_axi_out_V_ARADDR => open,
    m_axi_out_V_ARID => open,
    m_axi_out_V_ARLEN => open,
    m_axi_out_V_ARSIZE => open,
    m_axi_out_V_ARBURST => open,
    m_axi_out_V_ARLOCK => open,
    m_axi_out_V_ARCACHE => open,
    m_axi_out_V_ARPROT => open,
    m_axi_out_V_ARQOS => open,
    m_axi_out_V_ARREGION => open,
    m_axi_out_V_ARUSER => open,
    m_axi_out_V_RVALID => '0',
    m_axi_out_V_RREADY => open,
    m_axi_out_V_RDATA => ap_const_lv512_lc_1,
    m_axi_out_V_RLAST => '0',
    m_axi_out_V_RID => "0",
    m_axi_out_V_RUSER => "0",
    m_axi_out_V_RRESP => "00",
    m_axi_out_V_BVALID => write_output_m_axi_out_V_BVALID,
    m_axi_out_V_BREADY => write_output_m_axi_out_V_BREADY,
    m_axi_out_V_BRESP => write_output_m_axi_out_V_BRESP,
    m_axi_out_V_BID => write_output_m_axi_out_V_BID,
    m_axi_out_V_BUSER => write_output_m_axi_out_V_BUSER,
    out_V_offset => reg_mem_offset_shifted,
    address => reg_address,
    data_len => reg_data_len
  );

  -- AXI interface
  hls_m_axi_i: entity work.hls_sdaccel_kernel_iostreams_hls_gmem0_m_axi
  generic map (
    CONSERVATIVE => 0,
    USER_DW => 512,
    USER_AW => 64,
    USER_MAXREQS => 8,           -- do not set below 2
    NUM_READ_OUTSTANDING => 2,   -- do not set below 2 - no reads in this module
    NUM_WRITE_OUTSTANDING => 8,  -- do not set below 2
    MAX_READ_BURST_LENGTH => 2,  -- no reads in this module
    MAX_WRITE_BURST_LENGTH => 16,
    C_M_AXI_ID_WIDTH => C_M_AXI_GMEMWRITE_ID_WIDTH,
    C_M_AXI_ADDR_WIDTH => C_M_AXI_GMEMWRITE_ADDR_WIDTH,
    C_TARGET_ADDR => 16#00000000#,
    C_M_AXI_DATA_WIDTH => C_M_AXI_GMEMWRITE_DATA_WIDTH,
    C_M_AXI_AWUSER_WIDTH => C_M_AXI_GMEMWRITE_AWUSER_WIDTH,
    C_M_AXI_ARUSER_WIDTH => C_M_AXI_GMEMWRITE_ARUSER_WIDTH,
    C_M_AXI_WUSER_WIDTH => C_M_AXI_GMEMWRITE_WUSER_WIDTH,
    C_M_AXI_RUSER_WIDTH => C_M_AXI_GMEMWRITE_RUSER_WIDTH,
    C_M_AXI_BUSER_WIDTH => C_M_AXI_GMEMWRITE_BUSER_WIDTH,
    C_USER_VALUE => C_M_AXI_GMEMWRITE_USER_VALUE,
    C_PROT_VALUE => C_M_AXI_GMEMWRITE_PROT_VALUE,
    C_CACHE_VALUE => C_M_AXI_GMEMWRITE_CACHE_VALUE)
  port map (
    ACLK => clk_axi,
    ARESET => rst_axi,
    ACLK_EN => '1',
    AWVALID => m_axi_gmem_AWVALID,
    AWREADY => m_axi_gmem_AWREADY,
    AWADDR => m_axi_gmem_AWADDR,
    AWID => m_axi_gmem_AWID,
    AWLEN => m_axi_gmem_AWLEN,
    AWSIZE => m_axi_gmem_AWSIZE,
    AWBURST => m_axi_gmem_AWBURST,
    AWLOCK => m_axi_gmem_AWLOCK,
    AWCACHE => m_axi_gmem_AWCACHE,
    AWPROT => m_axi_gmem_AWPROT,
    AWQOS => m_axi_gmem_AWQOS,
    AWREGION => m_axi_gmem_AWREGION,
    AWUSER => m_axi_gmem_AWUSER,
    WVALID => m_axi_gmem_WVALID,
    WREADY => m_axi_gmem_WREADY,
    WDATA => m_axi_gmem_WDATA,
    WSTRB => m_axi_gmem_WSTRB,
    WLAST => m_axi_gmem_WLAST,
    WID => m_axi_gmem_WID,
    WUSER => m_axi_gmem_WUSER,
    ARVALID => m_axi_gmem_ARVALID,
    ARREADY => m_axi_gmem_ARREADY,
    ARADDR => m_axi_gmem_ARADDR,
    ARID => m_axi_gmem_ARID,
    ARLEN => m_axi_gmem_ARLEN,
    ARSIZE => m_axi_gmem_ARSIZE,
    ARBURST => m_axi_gmem_ARBURST,
    ARLOCK => m_axi_gmem_ARLOCK,
    ARCACHE => m_axi_gmem_ARCACHE,
    ARPROT => m_axi_gmem_ARPROT,
    ARQOS => m_axi_gmem_ARQOS,
    ARREGION => m_axi_gmem_ARREGION,
    ARUSER => m_axi_gmem_ARUSER,
    RVALID => m_axi_gmem_RVALID,
    RREADY => m_axi_gmem_RREADY,
    RDATA => m_axi_gmem_RDATA,
    RLAST => m_axi_gmem_RLAST,
    RID => m_axi_gmem_RID,
    RUSER => m_axi_gmem_RUSER,
    RRESP => m_axi_gmem_RRESP,
    BVALID => m_axi_gmem_BVALID,
    BREADY => m_axi_gmem_BREADY,
    BRESP => m_axi_gmem_BRESP,
    BID => m_axi_gmem_BID,
    BUSER => m_axi_gmem_BUSER,
    -- internal bus ports
    -- read channel is disabled for this module
    I_AWVALID => write_output_m_axi_out_V_AWVALID,
    I_AWREADY => write_output_m_axi_out_V_AWREADY,
    I_AWADDR => write_output_m_axi_out_V_AWADDR,
    I_AWID => write_output_m_axi_out_V_AWID,
    I_AWLEN => write_output_m_axi_out_V_AWLEN,
    I_AWSIZE => write_output_m_axi_out_V_AWSIZE,
    I_AWLOCK => write_output_m_axi_out_V_AWLOCK,
    I_AWCACHE => write_output_m_axi_out_V_AWCACHE,
    I_AWQOS => write_output_m_axi_out_V_AWQOS,
    I_AWPROT => write_output_m_axi_out_V_AWPROT,
    I_AWUSER => write_output_m_axi_out_V_AWUSER,
    I_AWBURST => write_output_m_axi_out_V_AWBURST,
    I_AWREGION => write_output_m_axi_out_V_AWREGION,
    I_WVALID => write_output_m_axi_out_V_WVALID,
    I_WREADY => write_output_m_axi_out_V_WREADY,
    I_WDATA => write_output_m_axi_out_V_WDATA,
    I_WID => write_output_m_axi_out_V_WID,
    I_WUSER => write_output_m_axi_out_V_WUSER,
    I_WLAST => write_output_m_axi_out_V_WLAST,
    I_WSTRB => write_output_m_axi_out_V_WSTRB,
    I_ARVALID => '0',
    I_ARREADY => open,
    I_ARADDR => x"0000000000000000",
    I_ARID => "0",
    I_ARLEN => x"00000000",
    I_ARSIZE => "000",
    I_ARLOCK => "00",
    I_ARCACHE => "0000",
    I_ARQOS => "0000",
    I_ARPROT => "000",
    I_ARUSER => "0",
    I_ARBURST => "00",
    I_ARREGION => "0000",
    I_RVALID => open,
    I_RREADY => '0',
    I_RDATA => open,
    I_RID => open,
    I_RUSER => open,
    I_RRESP => open,
    I_RLAST => open,
    I_BVALID => write_output_m_axi_out_V_BVALID,
    I_BREADY => write_output_m_axi_out_V_BREADY,
    I_BRESP => write_output_m_axi_out_V_BRESP,
    I_BID => write_output_m_axi_out_V_BID,
    I_BUSER => write_output_m_axi_out_V_BUSER
  );

end architecture;

