../output-impl-vhdl/dataflow_in_loop.vhd