../output-impl-vhdl/write_stream_proc.vhd