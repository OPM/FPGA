../output-impl-vhdl/fifo_w512_d512_A_x.vhd