../output-impl-vhdl/write_output.vhd