../output-impl-vhdl/read_input.vhd