../output-impl-vhdl/start_for_write_stream_proc_U0.vhd