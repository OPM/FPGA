../output-impl-vhdl/hls_sdaccel_kernel_iostreams_hls_gmem0_m_axi.vhd