--  Copyright 2020 Equinor ASA
--
--  This file is part of the Open Porous Media project (OPM).
--
--  OPM is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  OPM is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with OPM.  If not, see <http://www.gnu.org/licenses/>.

-- *******************************
-- top for AXI memory write module
-- *******************************
-- WARNING: this design is meant for a write port connected to DDR memory.
-- This design integrates:
-- * the write_output core generated by HLS
-- * the AXI master core generated by HLS
-- * a FIFO that includes the almost_full signal (generated by HLS and modified)
-- * registers for address, data_len, offset when ap_start is set (HLS
--   module does not properly register them!)

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
library work;
  use work.axi_io_common.all;

entity mem_write_top_ddr is
port (
  -- HLS interface
  ap_clk : in std_logic;
  ap_rst : in std_logic;
  ap_start : in std_logic;
  ap_done : out std_logic;
  ap_idle : out std_logic;
  ap_ready : out std_logic;
  -- parameters
  address : in std_logic_vector (63 downto 0);
  data_len : in std_logic_vector (31 downto 0);
  -- AXI interface
  mem_offset : in std_logic_vector (63 downto 0);
  m_axi_gmem_AWVALID : out std_logic;
  m_axi_gmem_AWREADY : in std_logic;
  m_axi_gmem_AWADDR : out std_logic_vector (C_M_AXI_GMEMWRITE_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_AWID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_AWLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_AWSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_AWCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_AWQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_AWUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_AWUSER_WIDTH-1 downto 0);
  m_axi_gmem_WVALID : out std_logic;
  m_axi_gmem_WREADY : in std_logic;
  m_axi_gmem_WDATA : out std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH-1 downto 0);
  m_axi_gmem_WSTRB : out std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH/8-1 downto 0);
  m_axi_gmem_WLAST : out std_logic;
  m_axi_gmem_WID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_WUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_WUSER_WIDTH-1 downto 0);
  m_axi_gmem_ARVALID : out std_logic;
  m_axi_gmem_ARREADY : in std_logic;
  m_axi_gmem_ARADDR : out std_logic_vector (C_M_AXI_GMEMWRITE_ADDR_WIDTH-1 downto 0);
  m_axi_gmem_ARID : out std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_ARLEN : out std_logic_vector (7 downto 0);
  m_axi_gmem_ARSIZE : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARBURST : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARLOCK : out std_logic_vector (1 downto 0);
  m_axi_gmem_ARCACHE : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARPROT : out std_logic_vector (2 downto 0);
  m_axi_gmem_ARQOS : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARREGION : out std_logic_vector (3 downto 0);
  m_axi_gmem_ARUSER : out std_logic_vector (C_M_AXI_GMEMWRITE_ARUSER_WIDTH-1 downto 0);
  m_axi_gmem_RVALID : in std_logic;
  m_axi_gmem_RREADY : out std_logic;
  m_axi_gmem_RDATA : in std_logic_vector (C_M_AXI_GMEMWRITE_DATA_WIDTH-1 downto 0);
  m_axi_gmem_RLAST : in std_logic;
  m_axi_gmem_RID : in std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_RUSER : in std_logic_vector (C_M_AXI_GMEMWRITE_RUSER_WIDTH-1 downto 0);
  m_axi_gmem_RRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BVALID : in std_logic;
  m_axi_gmem_BREADY : out std_logic;
  m_axi_gmem_BRESP : in std_logic_vector (1 downto 0);
  m_axi_gmem_BID : in std_logic_vector (C_M_AXI_GMEMWRITE_ID_WIDTH-1 downto 0);
  m_axi_gmem_BUSER : in std_logic_vector (C_M_AXI_GMEMWRITE_BUSER_WIDTH-1 downto 0);
  -- FIFO (stream) interface
  out_fifo_data : in std_logic_vector(C_FIFOWRITE_DATAIN_WIDTH-1 downto 0);
  out_fifo_full : out std_logic;
  out_fifo_almost_full : out std_logic;
  out_fifo_wr : in std_logic
);
end;

architecture behavioral of mem_write_top_ddr is
signal reg_ap_start, reg_ap_done, reg_ap_idle, reg_ap_ready: std_logic;
signal reg_address: std_logic_vector (63 downto 0);
signal reg_data_len: std_logic_vector (31 downto 0);
signal reg_mem_offset_shifted: std_logic_vector(57 downto 0);
signal write_output_fifo_data: std_logic_vector(C_FIFOWRITE_DATAOUT_WIDTH-1 downto 0);
signal write_output_fifo_empty_n, write_output_fifo_rd: std_logic;
signal write_output_m_axi_out_V_AWVALID: std_logic;
signal write_output_m_axi_out_V_AWREADY: std_logic;
signal write_output_m_axi_out_V_AWADDR: std_logic_vector (63 downto 0);
signal write_output_m_axi_out_V_AWID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_AWLEN: std_logic_vector (31 downto 0);
signal write_output_m_axi_out_V_AWSIZE: std_logic_vector (2 downto 0);
signal write_output_m_axi_out_V_AWLOCK: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_AWCACHE: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_AWQOS: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_AWPROT: std_logic_vector (2 downto 0);
signal write_output_m_axi_out_V_AWUSER: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_AWBURST: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_AWREGION: std_logic_vector (3 downto 0);
signal write_output_m_axi_out_V_WVALID: std_logic;
signal write_output_m_axi_out_V_WREADY: std_logic;
signal write_output_m_axi_out_V_WDATA: std_logic_vector (511 downto 0);
signal write_output_m_axi_out_V_WID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_WUSER: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_WLAST: std_logic;
signal write_output_m_axi_out_V_WSTRB: std_logic_vector (63 downto 0);
signal write_output_m_axi_out_V_BVALID: std_logic;
signal write_output_m_axi_out_V_BREADY: std_logic;
signal write_output_m_axi_out_V_BRESP: std_logic_vector (1 downto 0);
signal write_output_m_axi_out_V_BID: std_logic_vector (0 downto 0);
signal write_output_m_axi_out_V_BUSER: std_logic_vector (0 downto 0);
type control_t is (idle,running);
-- number of words contained by the FIFO
constant FIFO_WORDS: integer := 512;

begin

  -- process to resync the signals that must be registered to fix the wrong
  -- bevahior of write_output unit
  -- uses single-shot style for ap_done
  control_os_p: process(ap_clk, ap_start)
  variable state: control_t;
  variable vready: std_logic;
  begin
    if rising_edge(ap_clk) then
      if ap_rst = '1' then
        ap_done <= '0';
        ap_ready <= '0';
        vready := '0';
        reg_ap_start <= '0';
        state := idle;
      else
        case state is
          when idle =>
            -- wait until ap_start is set
            ap_done <= '0';
            ap_ready <= '0';
            vready := '0';
            reg_ap_start <= '0';
            if (ap_start = '1') then
              reg_ap_start <= '1';
              reg_address <= address;
              reg_data_len <= data_len;
              reg_mem_offset_shifted <= mem_offset(63 downto 6);
              state := running;
            end if;
          when running =>
            -- run the unit
            reg_ap_start <= '0';
            if (reg_ap_done = '1') then
              ap_done <= '1';
              ap_ready <= '1';
              vready := '1';
              state := idle;
            end if;
          when others =>
            state := idle;
        end case;
      end if;
    end if;
    if (ap_start = '1') or (vready = '1') or (state = running) then
      ap_idle <= '0';
    else
      ap_idle <= '1';
    end if;
  end process;

  -- process to resync the signals that must be registered to fix the wrong
  -- bevahior of write_output unit
  -- uses SDx/HLS style for ap_done (stays set until next start is given)
--  control_sdx_p: process(ap_clk, ap_start)
--  variable state: control_t;
--  variable vready: std_logic;
--  begin
--    if rising_edge(ap_clk) then
--      if ap_rst = '1' then
--        ap_ready <= '0';
--        vready := '0';
--        reg_ap_start <= '0';
--        state := idle;
--      else
--        case state is
--          when idle =>
--            -- wait until ap_start is set
--            ap_ready <= '0';
--            vready := '0';
--            reg_ap_start <= '0';
--            if (ap_start = '1') then
--              reg_ap_start <= '1';
--              reg_address <= address;
--              reg_data_len <= data_len;
--              reg_mem_offset_shifted <= mem_offset(63 downto 6);
--              state := running;
--            end if;
--          when running =>
--            -- run the unit
--            reg_ap_start <= '0';
--            if (reg_ap_done = '1') then
--              ap_ready <= '1';
--              vready := '1';
--              state := idle;
--            end if;
--          when others =>
--            state := idle;
--        end case;
--      end if;
--    end if;
--    if (ap_start = '1') or (state = running) then
--      ap_done <= '0';
--    else
--      ap_done <= '1';
--    end if;
--    if (ap_start = '1') or (vready = '1') or (state = running) then
--      ap_idle <= '0';
--    else
--      ap_idle <= '1';
--    end if;
--  end process;

  -- AXI interface
  hls_m_axi_i: entity work.hls_sdaccel_kernel_iostreams_hls_gmem0_m_axi
  generic map (
    CONSERVATIVE => 0,
    USER_DW => 512,
    USER_AW => 64,
    USER_MAXREQS => 8,           -- do not set below 2
    NUM_READ_OUTSTANDING => 2,   -- do not set below 2 - no reads in this module
    NUM_WRITE_OUTSTANDING => 8,  -- do not set below 2
    MAX_READ_BURST_LENGTH => 2,  -- no reads in this module
    MAX_WRITE_BURST_LENGTH => 256,
    C_M_AXI_ID_WIDTH => C_M_AXI_GMEMWRITE_ID_WIDTH,
    C_M_AXI_ADDR_WIDTH => C_M_AXI_GMEMWRITE_ADDR_WIDTH,
    C_TARGET_ADDR => 16#00000000#,
    C_M_AXI_DATA_WIDTH => C_M_AXI_GMEMWRITE_DATA_WIDTH,
    C_M_AXI_AWUSER_WIDTH => C_M_AXI_GMEMWRITE_AWUSER_WIDTH,
    C_M_AXI_ARUSER_WIDTH => C_M_AXI_GMEMWRITE_ARUSER_WIDTH,
    C_M_AXI_WUSER_WIDTH => C_M_AXI_GMEMWRITE_WUSER_WIDTH,
    C_M_AXI_RUSER_WIDTH => C_M_AXI_GMEMWRITE_RUSER_WIDTH,
    C_M_AXI_BUSER_WIDTH => C_M_AXI_GMEMWRITE_BUSER_WIDTH,
    C_USER_VALUE => C_M_AXI_GMEMWRITE_USER_VALUE,
    C_PROT_VALUE => C_M_AXI_GMEMWRITE_PROT_VALUE,
    C_CACHE_VALUE => C_M_AXI_GMEMWRITE_CACHE_VALUE)
  port map (
    ACLK => ap_clk,
    ARESET => ap_rst,
    ACLK_EN => '1',
    AWVALID => m_axi_gmem_AWVALID,
    AWREADY => m_axi_gmem_AWREADY,
    AWADDR => m_axi_gmem_AWADDR,
    AWID => m_axi_gmem_AWID,
    AWLEN => m_axi_gmem_AWLEN,
    AWSIZE => m_axi_gmem_AWSIZE,
    AWBURST => m_axi_gmem_AWBURST,
    AWLOCK => m_axi_gmem_AWLOCK,
    AWCACHE => m_axi_gmem_AWCACHE,
    AWPROT => m_axi_gmem_AWPROT,
    AWQOS => m_axi_gmem_AWQOS,
    AWREGION => m_axi_gmem_AWREGION,
    AWUSER => m_axi_gmem_AWUSER,
    WVALID => m_axi_gmem_WVALID,
    WREADY => m_axi_gmem_WREADY,
    WDATA => m_axi_gmem_WDATA,
    WSTRB => m_axi_gmem_WSTRB,
    WLAST => m_axi_gmem_WLAST,
    WID => m_axi_gmem_WID,
    WUSER => m_axi_gmem_WUSER,
    ARVALID => m_axi_gmem_ARVALID,
    ARREADY => m_axi_gmem_ARREADY,
    ARADDR => m_axi_gmem_ARADDR,
    ARID => m_axi_gmem_ARID,
    ARLEN => m_axi_gmem_ARLEN,
    ARSIZE => m_axi_gmem_ARSIZE,
    ARBURST => m_axi_gmem_ARBURST,
    ARLOCK => m_axi_gmem_ARLOCK,
    ARCACHE => m_axi_gmem_ARCACHE,
    ARPROT => m_axi_gmem_ARPROT,
    ARQOS => m_axi_gmem_ARQOS,
    ARREGION => m_axi_gmem_ARREGION,
    ARUSER => m_axi_gmem_ARUSER,
    RVALID => m_axi_gmem_RVALID,
    RREADY => m_axi_gmem_RREADY,
    RDATA => m_axi_gmem_RDATA,
    RLAST => m_axi_gmem_RLAST,
    RID => m_axi_gmem_RID,
    RUSER => m_axi_gmem_RUSER,
    RRESP => m_axi_gmem_RRESP,
    BVALID => m_axi_gmem_BVALID,
    BREADY => m_axi_gmem_BREADY,
    BRESP => m_axi_gmem_BRESP,
    BID => m_axi_gmem_BID,
    BUSER => m_axi_gmem_BUSER,
    -- internal bus ports
    -- read channel is disabled for this module
    I_AWVALID => write_output_m_axi_out_V_AWVALID,
    I_AWREADY => write_output_m_axi_out_V_AWREADY,
    I_AWADDR => write_output_m_axi_out_V_AWADDR,
    I_AWID => write_output_m_axi_out_V_AWID,
    I_AWLEN => write_output_m_axi_out_V_AWLEN,
    I_AWSIZE => write_output_m_axi_out_V_AWSIZE,
    I_AWLOCK => write_output_m_axi_out_V_AWLOCK,
    I_AWCACHE => write_output_m_axi_out_V_AWCACHE,
    I_AWQOS => write_output_m_axi_out_V_AWQOS,
    I_AWPROT => write_output_m_axi_out_V_AWPROT,
    I_AWUSER => write_output_m_axi_out_V_AWUSER,
    I_AWBURST => write_output_m_axi_out_V_AWBURST,
    I_AWREGION => write_output_m_axi_out_V_AWREGION,
    I_WVALID => write_output_m_axi_out_V_WVALID,
    I_WREADY => write_output_m_axi_out_V_WREADY,
    I_WDATA => write_output_m_axi_out_V_WDATA,
    I_WID => write_output_m_axi_out_V_WID,
    I_WUSER => write_output_m_axi_out_V_WUSER,
    I_WLAST => write_output_m_axi_out_V_WLAST,
    I_WSTRB => write_output_m_axi_out_V_WSTRB,
    I_ARVALID => '0',
    I_ARREADY => open,
    I_ARADDR => x"0000000000000000",
    I_ARID => "0",
    I_ARLEN => x"00000000",
    I_ARSIZE => "000",
    I_ARLOCK => "00",
    I_ARCACHE => "0000",
    I_ARQOS => "0000",
    I_ARPROT => "000",
    I_ARUSER => "0",
    I_ARBURST => "00",
    I_ARREGION => "0000",
    I_RVALID => open,
    I_RREADY => '0',
    I_RDATA => open,
    I_RID => open,
    I_RUSER => open,
    I_RRESP => open,
    I_RLAST => open,
    I_BVALID => write_output_m_axi_out_V_BVALID,
    I_BREADY => write_output_m_axi_out_V_BREADY,
    I_BRESP => write_output_m_axi_out_V_BRESP,
    I_BID => write_output_m_axi_out_V_BID,
    I_BUSER => write_output_m_axi_out_V_BUSER
  );

  -- memory write module
  write_output_i: entity work.write_output
  port map (
    ap_clk => ap_clk,
    ap_rst => ap_rst,
    ap_start => reg_ap_start,
    ap_done => reg_ap_done,
    ap_idle => reg_ap_idle,
    ap_ready => reg_ap_ready,
    resultStream_V_V_dout => write_output_fifo_data,
    resultStream_V_V_empty_n => write_output_fifo_empty_n,
    resultStream_V_V_read => write_output_fifo_rd,
    m_axi_out_V_AWVALID => write_output_m_axi_out_V_AWVALID,
    m_axi_out_V_AWREADY => write_output_m_axi_out_V_AWREADY,
    m_axi_out_V_AWADDR => write_output_m_axi_out_V_AWADDR,
    m_axi_out_V_AWID => write_output_m_axi_out_V_AWID,
    m_axi_out_V_AWLEN => write_output_m_axi_out_V_AWLEN,
    m_axi_out_V_AWSIZE => write_output_m_axi_out_V_AWSIZE,
    m_axi_out_V_AWBURST => write_output_m_axi_out_V_AWBURST,
    m_axi_out_V_AWLOCK => write_output_m_axi_out_V_AWLOCK,
    m_axi_out_V_AWCACHE => write_output_m_axi_out_V_AWCACHE,
    m_axi_out_V_AWPROT => write_output_m_axi_out_V_AWPROT,
    m_axi_out_V_AWQOS => write_output_m_axi_out_V_AWQOS,
    m_axi_out_V_AWREGION => write_output_m_axi_out_V_AWREGION,
    m_axi_out_V_AWUSER => write_output_m_axi_out_V_AWUSER,
    m_axi_out_V_WVALID => write_output_m_axi_out_V_WVALID,
    m_axi_out_V_WREADY => write_output_m_axi_out_V_WREADY,
    m_axi_out_V_WDATA => write_output_m_axi_out_V_WDATA,
    m_axi_out_V_WSTRB => write_output_m_axi_out_V_WSTRB,
    m_axi_out_V_WLAST => write_output_m_axi_out_V_WLAST,
    m_axi_out_V_WID => write_output_m_axi_out_V_WID,
    m_axi_out_V_WUSER => write_output_m_axi_out_V_WUSER,
    m_axi_out_V_ARVALID => open,
    m_axi_out_V_ARREADY => '0',
    m_axi_out_V_ARADDR => open,
    m_axi_out_V_ARID => open,
    m_axi_out_V_ARLEN => open,
    m_axi_out_V_ARSIZE => open,
    m_axi_out_V_ARBURST => open,
    m_axi_out_V_ARLOCK => open,
    m_axi_out_V_ARCACHE => open,
    m_axi_out_V_ARPROT => open,
    m_axi_out_V_ARQOS => open,
    m_axi_out_V_ARREGION => open,
    m_axi_out_V_ARUSER => open,
    m_axi_out_V_RVALID => '0',
    m_axi_out_V_RREADY => open,
    m_axi_out_V_RDATA => ap_const_lv512_lc_1,
    m_axi_out_V_RLAST => '0',
    m_axi_out_V_RID => "0",
    m_axi_out_V_RUSER => "0",
    m_axi_out_V_RRESP => "00",
    m_axi_out_V_BVALID => write_output_m_axi_out_V_BVALID,
    m_axi_out_V_BREADY => write_output_m_axi_out_V_BREADY,
    m_axi_out_V_BRESP => write_output_m_axi_out_V_BRESP,
    m_axi_out_V_BID => write_output_m_axi_out_V_BID,
    m_axi_out_V_BUSER => write_output_m_axi_out_V_BUSER,
    out_V_offset => reg_mem_offset_shifted,
    address => reg_address,
    data_len => reg_data_len
  );

  -- write data FIFO
  outdata_fifo_i: entity work.fifo_out_w512
  generic map (
    MEM_STYLE  => "block",
    DATA_WIDTH => 512,
    DEPTH      => FIFO_WORDS)
  port map (
    clk => ap_clk,
    reset => ap_rst,
    if_almost_full => out_fifo_almost_full,
    if_full => out_fifo_full,
    if_write_ce => '1',
    if_write => out_fifo_wr,
    if_din => out_fifo_data,
    if_empty_n => write_output_fifo_empty_n,
    if_read_ce => '1',
    if_read => write_output_fifo_rd,
    if_dout => write_output_fifo_data
  );

end architecture;

