../output-impl-vhdl/fifo_w10_d2_A.vhd